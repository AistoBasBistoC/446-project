`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/06/2021 05:42:58 AM
// Design Name: 
// Module Name: Top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Top(
    input Clk, Reset,
    input [7:0] AN,
    output [7:0] display,
    output [7:0] Anode
    );
    
    
    assign Anode = AN;
    /// Connect different building block together
	
	wire Clock1Hz;
    wire [3:0] Count;
    
    assign Anode = AN;
    /// Connect different building block together
    
    //1. Clock Divider 1Hz Frequency
    Clock_Divider BLOCK1 (.Clk(Clk), .Reset(Reset), .Slow_Clock(Clock1Hz));
    
    //2. Counter 0-9
    //Counter is driven by  slow clock generated by clock divider 
    Counter BLOCK2 (.Clk(Clock1Hz), .Reset(Reset),.Q(Count));
    
    //3. Binary to 7 segment
    Bin_7Segment BLOCK3 (.Bin(Count), .Seven_Segment(display));
    
endmodule
