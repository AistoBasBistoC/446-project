`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/06/2021 05:36:58 AM
// Design Name: 
// Module Name: Counter
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Counter(
    input Clk, Reset,
    output [3:0] Q
    );
    
// Make sure your Counter is driven by  slow clock generated by clock divider
parameter ST_ZERO = 4’b0000, ST_ONE = 4’b0001, ST_TWO = 4’b0010, ST_THREE = 4’b0011, ST_FOUR = 4’b0100, ST_FIVE = 4’b0101, ST_SIX = 4’b0110, ST_SEVEN = 4’b0111, ST_EIGHT = 4’b1000, ST_NINE = 4’b1001;

reg [3:0] state, n_state; //state = present state, n_state = next state

always @(posedge Clk, posedge Reset)
	if (Reset)
		state <= ST_ZERO;
		else
		state <= n_state;

always @(*)
	case (state)
		ST_ZERO: 
			n_state <= ST_ONE;			
		ST_ONE: 
			n_state <= ST_TWO;
		ST_TWO: 
			n_state <= ST_THREE;
		ST_THREE: 
			n_state <= ST_FOUR;
		ST_FOUR: 
			n_state <= ST_FIVE;
		ST_FIVE: 
			n_state <= ST_SIX;
		ST_SIX: 
			n_state <= ST_SEVEN;
		ST_SEVEN: 
			n_state <= ST_EIGHT;
		ST_EIGHT: 
			n_state <= ST_NINE;
		ST_NINE: 
			n_state <= ST_ZERO;
		default: 
			n_state <= ST_ZERO;
	endcase

assign Q = state;

endmodule

