`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/06/2021 05:36:58 AM
// Design Name: 
// Module Name: Counter
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Counter(
    input Clk, Reset,
    output [3:0] Q
    );
    
    // Make sure your Counter is driven by  slow clock generated by clock divider
    always @(posedge Clk) begin 
	if (!Reset)
		Q <= 1’b0;
	else
		Q <= Q + 1’b1;
end  
endmodule
