`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/06/2021 05:36:58 AM
// Design Name: 
// Module Name: Counter
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Counter(
    input Clk, Reset,
    output [3:0] Q
    );
    reg [3:0] PS, NS;   //PS = Present State, NS = Next State
    
    // Make sure your Counter is driven by  slow clock generated by clock divider
    
    //state declarations
    parameter S0 = 4'b0000; //0
    parameter S1 = 4'b0001; //1
    parameter S2 = 4'b0010; //2
    parameter S3 = 4'b0011; //3
    parameter S4 = 4'b0100; //4
    parameter S5 = 4'b0101; //5
    parameter S6 = 4'b0110; //6
    parameter S7 = 4'b0111; //7
    parameter S8 = 4'b1000; //8
    parameter S9 = 4'b1001; //9
    
    //Reset Check
    always @(posedge Clk, posedge Reset)
        if(Reset) PS <= S0;
        else
        PS <= NS;
        
    //Machine State Transitions
    always@(*)
    case(PS)
    S0: NS = S1;
    S1: NS = S2;
    S2: NS = S3;
    S3: NS = S4;
    S4: NS = S5;
    S5: NS = S6;
    S6: NS = S7;
    S7: NS = S8;
    S8: NS = S9;
    S9: NS = S0;
    default: NS = S0;
    endcase
    
    assign Q = PS;
    
endmodule
