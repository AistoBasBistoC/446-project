`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/06/2021 05:36:58 AM
// Design Name: 
// Module Name: Counter
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Counter(
    input Clk, Reset,
    output [3:0] Q
    );
    
// Make sure your Counter is driven by  slow clock generated by clock divider
parameter ST_ZERO = 4’b0000, ST_ONE = 4’b0001, ST_TWO = 4’b0010, ST_THREE = 4’b0011, ST_FOUR = 4’b0100, ST_FIVE = 4’b0101, ST_SIX = 4’b0110, ST_SEVEN = 4’b0111, ST_EIGHT = 4’b1000, ST_NINE = 4’b1001;

reg [3:0] state;

always @(posedge Clk or posedge Reset)
begin
	if (Reset == 1’b1) begin
		state = ST_ZERO;
		Q = 4’b0000;
	end else begin
	case (state)
		ST_ZERO: begin
			state = ST_ONE;
			Q = 4’b0000;
			end
		ST_ONE: begin
			state = ST_TWO;
			Q = 4’b0001;
			end
		ST_TWO: begin
			state = ST_THREE;
			Q = 4’b0010;
			end
		ST_THREE: begin
			state = ST_FOUR;
			Q = 4’b0011;
			end
		ST_FOUR: begin
			state = ST_FIVE;
			Q = 4’b0100;
			end
		ST_FIVE: begin
			state = ST_SIX;
			Q = 4’b0101;
			end
		ST_SIX: begin
			state = ST_SEVEN;
			Q = 4’b0110;
			end
		ST_SEVEN: begin
			state = ST_EIGHT;
			Q = 4’b0111;
			end
		ST_EIGHT: begin
			state = ST_NINE;
			Q = 4’b1000;
			end
		ST_NINE: begin
			state = ST_ZERO;
			Q = 4’b1001;
		default: begin
			state = ST_ZERO;
			Q = 4’b0000;
			end
		endcase
	end
end
endmodule

